`include "Async_fifo_memory.sv"
`include "rempty.sv"
`include "sync_rtow_wtor.sv"
`include "Wfull.sv"
`include "Fifo_top.sv"