package data_fields;

parameter DATASIZE=8;

endpackage